`timescale 1ns / 1ps
module kr260_top(
    output led
    );
    
    assign led = 1'b1;
    
endmodule
